/**
 * This file is part of the Coyote <https://github.com/fpgasystems/Coyote>
 *
 * MIT Licence
 * Copyright (c) 2025-2026, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

// Simple pipeline stages, buffering the input/output signals (not really needed, but nice to have for easier timing closure)
AXI4SR axis_in_int (.*);
axisr_reg inst_reg_in  (.aclk(aclk), .aresetn(aresetn), .s_axis(axis_host_recv[0]), .m_axis(axis_in_int));

AXI4SR axis_out_int (.*);
axisr_reg inst_reg_out (.aclk(aclk), .aresetn(aresetn), .s_axis(axis_out_int), .m_axis(axis_host_send[0]));

///////////////////////////////////////
//          BENCH CONTROL           //
/////////////////////////////////////
// Starting read/write operations
logic [1:0] bench_ctrl;
parameter integer START_RD = 0;
parameter integer START_WR = 1;

///////////////////////////////////////
//       COMMAND COMPLETION         //
/////////////////////////////////////
// Number of requested reads/writes; controlled by the user from software
// e.g., for latency we might do 1 and for throughput we might do 32
logic [31:0] bench_n_reps;

// Number of issued reads/writes
logic [31:0] bench_sent;

// Asserted high when all the commands have been marked as completed
logic done_req;

///////////////////////////////////////
//         DATA COMPLETION          //
/////////////////////////////////////
// Number of incoming/outgoing AXI data streams; 
// e.g. for a message of size 4096 bytes, the valid from the AXI stream goes high eight times
// and for 32 transfers (bench_n_reps = 32) like that, there will be 256 beats
// Set from the software to avoid computing divsion on the FPGA
logic [63:0] bench_n_beats;

// Number of completed AXI beats
logic [63:0] cnt_data;

// Asserted high when all the data has been processed
logic done_data;

///////////////////////////////////////
//        READ/WRITE DATA           //
/////////////////////////////////////
// Buffer size in bytes
logic [LEN_BITS-1:0] bench_len;

// Virtual address of buffer to be read from / written to
logic [VADDR_BITS-1:0] bench_vaddr;

// Coyote thread ID (obtained in software from coyote_thread.getCtid())
logic [PID_BITS-1:0] bench_pid;

///////////////////////////////////////
//           FSM & TIMING           //
/////////////////////////////////////
// In this example, reads and writes are de-coupled;
// That is, we either read bench_n_reps time from the buffer at bench_vaddr of size bench_len
// OR we write to the buffer of size bench_len at bench_vaddr; bench_n_reps times 
logic [1:0] state_C;
typedef enum logic[1:0]  {ST_IDLE, ST_READ, ST_WRITE} state_t;

// The values above are set from the software and propagated to the FPGA via PCIe and XDMA in a AXI Lite interface
// The helper module parses the AXI interface to the target signals
perf_fpga_axi_ctrl_parser inst_axi_ctrl_parser (
    .aclk(aclk),
    .aresetn(aresetn),
    .axi_ctrl(axi_ctrl),
    .bench_ctrl(bench_ctrl),
    .bench_pid(bench_pid),
    .bench_vaddr(bench_vaddr),
    .bench_len(bench_len),
    .bench_n_reps(bench_n_reps),
    .bench_n_beats(bench_n_beats)
);

// State-machine transition and counters
always_ff @(posedge aclk) begin
    if(aresetn == 1'b0) begin
        state_C <= ST_IDLE;
        cnt_data <= 0;
        bench_sent <= 0;

        done_req <= 1'b0;
        done_data <= 1'b0;

    end else begin
        case(state_C) 
            ST_IDLE: begin
                // Transition to next state if user triggered benchmark start
                state_C <= bench_ctrl[START_RD] ? ST_READ : 
                           bench_ctrl[START_WR] ? ST_WRITE : ST_IDLE;

                // Reset signals for new benchmark
                cnt_data <= 0;
                bench_sent <= 0;

                done_req <= 1'b0;
                done_data <= 1'b0;
            end
            ST_READ: begin
                // Request counter and completion
                bench_sent <= (sq_rd.valid && sq_rd.ready) ? bench_sent + 1 : bench_sent;
                done_req <= ((bench_sent == bench_n_reps - 1) && sq_rd.ready) ? 1'b1 : done_req;

                // Data counter and completion
                cnt_data <= (axis_in_int.tvalid && axis_in_int.tready) ? cnt_data + 1 : cnt_data;
                done_data <= ((cnt_data == bench_n_beats - 1) && axis_in_int.tvalid) ? 1'b1 : done_data;

                // Transition back to IDLE if complete; otherwise continue reading
                state_C <= (done_req && done_data) ? ST_IDLE : ST_READ;
            end
            ST_WRITE: begin
                // Request counter and completion
                done_req <= ((bench_sent == bench_n_reps - 1) && sq_wr.ready) ? 1'b1 : done_req;
                bench_sent <= (sq_wr.valid && sq_wr.ready) ? bench_sent + 1 : bench_sent;

                // Data counter and completion
                cnt_data <= (axis_out_int.tvalid && axis_out_int.tready) ? cnt_data + 1 : cnt_data;
                done_data <= ((cnt_data == bench_n_beats - 1) && axis_out_int.tready) ? 1'b1 : done_data;

                // Transition back to IDLE if complete; otherwise continue writing
                state_C <= (done_req && done_data) ? ST_IDLE : ST_WRITE;
            end
        endcase
    end
end

always_comb begin
    ///////////////////////////////
    //          READS           //
    /////////////////////////////
    // Requests
    sq_rd.data = 0;
    sq_rd.data.last = bench_sent == bench_n_reps - 1;
    sq_rd.data.pid = bench_pid;
    sq_rd.data.len = bench_len;
    sq_rd.data.vaddr = bench_vaddr;
    sq_rd.data.strm = STRM_HOST;
    sq_rd.data.opcode = LOCAL_READ;
    sq_rd.valid = (state_C == ST_READ) && ~done_req;

    cq_rd.ready = 1'b1;

    // Data
    axis_in_int.tready = (state_C == ST_READ) && ~done_data;

    ///////////////////////////////
    //          WRITES          //
    /////////////////////////////
    // Requests
    sq_wr.data = 0;
    sq_wr.data.last = bench_sent == bench_n_reps - 1;
    sq_wr.data.pid = bench_pid;
    sq_wr.data.len = bench_len;
    sq_wr.data.vaddr = bench_vaddr;
    sq_wr.data.strm = STRM_HOST;
    sq_wr.data.opcode = LOCAL_WRITE;
    sq_wr.valid = (state_C == ST_WRITE) && ~done_req;

    cq_wr.ready = 1'b1;

    // Data
    axis_out_int.tdata = cnt_data + 1;
    axis_out_int.tkeep = ~0;
    axis_out_int.tid   = 0;
    axis_out_int.tlast = cnt_data == bench_n_beats - 1;
    axis_out_int.tvalid = (state_C == ST_WRITE) && ~done_data;
end

// Tie off unused interfaces
always_comb notify.tie_off_m();
